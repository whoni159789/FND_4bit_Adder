`timescale 1ns / 1ps

module tb_BCD_TO_FND_Decoder();

    input i_EN;
    input [3:0] i_Value;
    output [7:0] o_Font;

    
endmodule
